-- multicore.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity multicore is
	port (
		clk_clk                     : in    std_logic                     := '0';             --                   clk.clk
		reset_reset_n               : in    std_logic                     := '0';             --                 reset.reset_n
		sdram_clk_clk               : out   std_logic;                                        --             sdram_clk.clk
		sdram_controller_wire_addr  : out   std_logic_vector(12 downto 0);                    -- sdram_controller_wire.addr
		sdram_controller_wire_ba    : out   std_logic_vector(1 downto 0);                     --                      .ba
		sdram_controller_wire_cas_n : out   std_logic;                                        --                      .cas_n
		sdram_controller_wire_cke   : out   std_logic;                                        --                      .cke
		sdram_controller_wire_cs_n  : out   std_logic;                                        --                      .cs_n
		sdram_controller_wire_dq    : inout std_logic_vector(15 downto 0) := (others => '0'); --                      .dq
		sdram_controller_wire_dqm   : out   std_logic_vector(1 downto 0);                     --                      .dqm
		sdram_controller_wire_ras_n : out   std_logic;                                        --                      .ras_n
		sdram_controller_wire_we_n  : out   std_logic                                         --                      .we_n
	);
end entity multicore;

architecture rtl of multicore is
	component multicore_cpu_1 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component multicore_cpu_1;

	component multicore_cpu_2 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component multicore_cpu_2;

	component multicore_cpu_3 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component multicore_cpu_3;

	component multicore_cpu_4 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component multicore_cpu_4;

	component multicore_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component multicore_jtag_uart;

	component multicore_mutex is
		port (
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			clk           : in  std_logic                     := 'X';             -- clk
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			data_from_cpu : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read          : in  std_logic                     := 'X';             -- read
			write         : in  std_logic                     := 'X';             -- write
			data_to_cpu   : out std_logic_vector(31 downto 0);                    -- readdata
			address       : in  std_logic                     := 'X'              -- address
		);
	end component multicore_mutex;

	component multicore_onchip_memory2_0 is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component multicore_onchip_memory2_0;

	component multicore_performance_counter is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component multicore_performance_counter;

	component multicore_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component multicore_pll;

	component multicore_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component multicore_sdram_controller;

	component multicore_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component multicore_sysid;

	component multicore_timer1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component multicore_timer1;

	component multicore_mm_interconnect_0 is
		port (
			pll_outclk0_clk                                 : in  std_logic                     := 'X';             -- clk
			cpu_1_reset_reset_bridge_in_reset_reset         : in  std_logic                     := 'X';             -- reset
			cpu_1_data_master_address                       : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_1_data_master_waitrequest                   : out std_logic;                                        -- waitrequest
			cpu_1_data_master_byteenable                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_1_data_master_read                          : in  std_logic                     := 'X';             -- read
			cpu_1_data_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_1_data_master_readdatavalid                 : out std_logic;                                        -- readdatavalid
			cpu_1_data_master_write                         : in  std_logic                     := 'X';             -- write
			cpu_1_data_master_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_1_data_master_debugaccess                   : in  std_logic                     := 'X';             -- debugaccess
			cpu_1_instruction_master_address                : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_1_instruction_master_waitrequest            : out std_logic;                                        -- waitrequest
			cpu_1_instruction_master_read                   : in  std_logic                     := 'X';             -- read
			cpu_1_instruction_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_1_instruction_master_readdatavalid          : out std_logic;                                        -- readdatavalid
			cpu_2_data_master_address                       : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_2_data_master_waitrequest                   : out std_logic;                                        -- waitrequest
			cpu_2_data_master_byteenable                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_2_data_master_read                          : in  std_logic                     := 'X';             -- read
			cpu_2_data_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_2_data_master_readdatavalid                 : out std_logic;                                        -- readdatavalid
			cpu_2_data_master_write                         : in  std_logic                     := 'X';             -- write
			cpu_2_data_master_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_2_data_master_debugaccess                   : in  std_logic                     := 'X';             -- debugaccess
			cpu_2_instruction_master_address                : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_2_instruction_master_waitrequest            : out std_logic;                                        -- waitrequest
			cpu_2_instruction_master_read                   : in  std_logic                     := 'X';             -- read
			cpu_2_instruction_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_2_instruction_master_readdatavalid          : out std_logic;                                        -- readdatavalid
			cpu_3_data_master_address                       : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_3_data_master_waitrequest                   : out std_logic;                                        -- waitrequest
			cpu_3_data_master_byteenable                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_3_data_master_read                          : in  std_logic                     := 'X';             -- read
			cpu_3_data_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_3_data_master_readdatavalid                 : out std_logic;                                        -- readdatavalid
			cpu_3_data_master_write                         : in  std_logic                     := 'X';             -- write
			cpu_3_data_master_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_3_data_master_debugaccess                   : in  std_logic                     := 'X';             -- debugaccess
			cpu_3_instruction_master_address                : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_3_instruction_master_waitrequest            : out std_logic;                                        -- waitrequest
			cpu_3_instruction_master_read                   : in  std_logic                     := 'X';             -- read
			cpu_3_instruction_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_3_instruction_master_readdatavalid          : out std_logic;                                        -- readdatavalid
			cpu_4_data_master_address                       : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_4_data_master_waitrequest                   : out std_logic;                                        -- waitrequest
			cpu_4_data_master_byteenable                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_4_data_master_read                          : in  std_logic                     := 'X';             -- read
			cpu_4_data_master_readdata                      : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_4_data_master_readdatavalid                 : out std_logic;                                        -- readdatavalid
			cpu_4_data_master_write                         : in  std_logic                     := 'X';             -- write
			cpu_4_data_master_writedata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_4_data_master_debugaccess                   : in  std_logic                     := 'X';             -- debugaccess
			cpu_4_instruction_master_address                : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_4_instruction_master_waitrequest            : out std_logic;                                        -- waitrequest
			cpu_4_instruction_master_read                   : in  std_logic                     := 'X';             -- read
			cpu_4_instruction_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_4_instruction_master_readdatavalid          : out std_logic;                                        -- readdatavalid
			cpu_1_debug_mem_slave_address                   : out std_logic_vector(8 downto 0);                     -- address
			cpu_1_debug_mem_slave_write                     : out std_logic;                                        -- write
			cpu_1_debug_mem_slave_read                      : out std_logic;                                        -- read
			cpu_1_debug_mem_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_1_debug_mem_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_1_debug_mem_slave_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_1_debug_mem_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			cpu_1_debug_mem_slave_debugaccess               : out std_logic;                                        -- debugaccess
			cpu_2_debug_mem_slave_address                   : out std_logic_vector(8 downto 0);                     -- address
			cpu_2_debug_mem_slave_write                     : out std_logic;                                        -- write
			cpu_2_debug_mem_slave_read                      : out std_logic;                                        -- read
			cpu_2_debug_mem_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_2_debug_mem_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_2_debug_mem_slave_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_2_debug_mem_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			cpu_2_debug_mem_slave_debugaccess               : out std_logic;                                        -- debugaccess
			cpu_3_debug_mem_slave_address                   : out std_logic_vector(8 downto 0);                     -- address
			cpu_3_debug_mem_slave_write                     : out std_logic;                                        -- write
			cpu_3_debug_mem_slave_read                      : out std_logic;                                        -- read
			cpu_3_debug_mem_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_3_debug_mem_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_3_debug_mem_slave_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_3_debug_mem_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			cpu_3_debug_mem_slave_debugaccess               : out std_logic;                                        -- debugaccess
			cpu_4_debug_mem_slave_address                   : out std_logic_vector(8 downto 0);                     -- address
			cpu_4_debug_mem_slave_write                     : out std_logic;                                        -- write
			cpu_4_debug_mem_slave_read                      : out std_logic;                                        -- read
			cpu_4_debug_mem_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_4_debug_mem_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_4_debug_mem_slave_byteenable                : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_4_debug_mem_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			cpu_4_debug_mem_slave_debugaccess               : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write               : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect          : out std_logic;                                        -- chipselect
			mutex_s1_address                                : out std_logic_vector(0 downto 0);                     -- address
			mutex_s1_write                                  : out std_logic;                                        -- write
			mutex_s1_read                                   : out std_logic;                                        -- read
			mutex_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mutex_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			mutex_s1_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_address                     : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory2_0_s1_write                       : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                  : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                       : out std_logic;                                        -- clken
			onchip_memory2_0_s2_address                     : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory2_0_s2_write                       : out std_logic;                                        -- write
			onchip_memory2_0_s2_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s2_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s2_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s2_chipselect                  : out std_logic;                                        -- chipselect
			onchip_memory2_0_s2_clken                       : out std_logic;                                        -- clken
			performance_counter_control_slave_address       : out std_logic_vector(3 downto 0);                     -- address
			performance_counter_control_slave_write         : out std_logic;                                        -- write
			performance_counter_control_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			performance_counter_control_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			performance_counter_control_slave_begintransfer : out std_logic;                                        -- begintransfer
			sdram_controller_s1_address                     : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                       : out std_logic;                                        -- write
			sdram_controller_s1_read                        : out std_logic;                                        -- read
			sdram_controller_s1_readdata                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                   : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                  : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid               : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                 : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                  : out std_logic;                                        -- chipselect
			sysid_control_slave_address                     : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer1_s1_address                               : out std_logic_vector(2 downto 0);                     -- address
			timer1_s1_write                                 : out std_logic;                                        -- write
			timer1_s1_readdata                              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer1_s1_writedata                             : out std_logic_vector(15 downto 0);                    -- writedata
			timer1_s1_chipselect                            : out std_logic;                                        -- chipselect
			timer_2_s1_address                              : out std_logic_vector(2 downto 0);                     -- address
			timer_2_s1_write                                : out std_logic;                                        -- write
			timer_2_s1_readdata                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_2_s1_writedata                            : out std_logic_vector(15 downto 0);                    -- writedata
			timer_2_s1_chipselect                           : out std_logic;                                        -- chipselect
			timer_3_s1_address                              : out std_logic_vector(2 downto 0);                     -- address
			timer_3_s1_write                                : out std_logic;                                        -- write
			timer_3_s1_readdata                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_3_s1_writedata                            : out std_logic_vector(15 downto 0);                    -- writedata
			timer_3_s1_chipselect                           : out std_logic;                                        -- chipselect
			timer_4_s1_address                              : out std_logic_vector(2 downto 0);                     -- address
			timer_4_s1_write                                : out std_logic;                                        -- write
			timer_4_s1_readdata                             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_4_s1_writedata                            : out std_logic_vector(15 downto 0);                    -- writedata
			timer_4_s1_chipselect                           : out std_logic                                         -- chipselect
		);
	end component multicore_mm_interconnect_0;

	component multicore_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component multicore_irq_mapper;

	component multicore_irq_mapper_001 is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component multicore_irq_mapper_001;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal pll_outclk0_clk                                                   : std_logic;                     -- pll:outclk_0 -> [cpu_1:clk, cpu_2:clk, cpu_3:clk, cpu_4:clk, irq_mapper:clk, irq_mapper_001:clk, irq_mapper_002:clk, irq_mapper_003:clk, jtag_uart:clk, mm_interconnect_0:pll_outclk0_clk, mutex:clk, onchip_memory2_0:clk, onchip_memory2_0:clk2, performance_counter:clk, rst_controller:clk, sdram_controller:clk, sysid:clock, timer1:clk, timer_2:clk, timer_3:clk, timer_4:clk]
	signal cpu_1_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_data_master_readdata -> cpu_1:d_readdata
	signal cpu_1_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_1_data_master_waitrequest -> cpu_1:d_waitrequest
	signal cpu_1_data_master_debugaccess                                     : std_logic;                     -- cpu_1:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_1_data_master_debugaccess
	signal cpu_1_data_master_address                                         : std_logic_vector(26 downto 0); -- cpu_1:d_address -> mm_interconnect_0:cpu_1_data_master_address
	signal cpu_1_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- cpu_1:d_byteenable -> mm_interconnect_0:cpu_1_data_master_byteenable
	signal cpu_1_data_master_read                                            : std_logic;                     -- cpu_1:d_read -> mm_interconnect_0:cpu_1_data_master_read
	signal cpu_1_data_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:cpu_1_data_master_readdatavalid -> cpu_1:d_readdatavalid
	signal cpu_1_data_master_write                                           : std_logic;                     -- cpu_1:d_write -> mm_interconnect_0:cpu_1_data_master_write
	signal cpu_1_data_master_writedata                                       : std_logic_vector(31 downto 0); -- cpu_1:d_writedata -> mm_interconnect_0:cpu_1_data_master_writedata
	signal cpu_2_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_2_data_master_readdata -> cpu_2:d_readdata
	signal cpu_2_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_2_data_master_waitrequest -> cpu_2:d_waitrequest
	signal cpu_2_data_master_debugaccess                                     : std_logic;                     -- cpu_2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_2_data_master_debugaccess
	signal cpu_2_data_master_address                                         : std_logic_vector(26 downto 0); -- cpu_2:d_address -> mm_interconnect_0:cpu_2_data_master_address
	signal cpu_2_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- cpu_2:d_byteenable -> mm_interconnect_0:cpu_2_data_master_byteenable
	signal cpu_2_data_master_read                                            : std_logic;                     -- cpu_2:d_read -> mm_interconnect_0:cpu_2_data_master_read
	signal cpu_2_data_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:cpu_2_data_master_readdatavalid -> cpu_2:d_readdatavalid
	signal cpu_2_data_master_write                                           : std_logic;                     -- cpu_2:d_write -> mm_interconnect_0:cpu_2_data_master_write
	signal cpu_2_data_master_writedata                                       : std_logic_vector(31 downto 0); -- cpu_2:d_writedata -> mm_interconnect_0:cpu_2_data_master_writedata
	signal cpu_3_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_3_data_master_readdata -> cpu_3:d_readdata
	signal cpu_3_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_3_data_master_waitrequest -> cpu_3:d_waitrequest
	signal cpu_3_data_master_debugaccess                                     : std_logic;                     -- cpu_3:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_3_data_master_debugaccess
	signal cpu_3_data_master_address                                         : std_logic_vector(26 downto 0); -- cpu_3:d_address -> mm_interconnect_0:cpu_3_data_master_address
	signal cpu_3_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- cpu_3:d_byteenable -> mm_interconnect_0:cpu_3_data_master_byteenable
	signal cpu_3_data_master_read                                            : std_logic;                     -- cpu_3:d_read -> mm_interconnect_0:cpu_3_data_master_read
	signal cpu_3_data_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:cpu_3_data_master_readdatavalid -> cpu_3:d_readdatavalid
	signal cpu_3_data_master_write                                           : std_logic;                     -- cpu_3:d_write -> mm_interconnect_0:cpu_3_data_master_write
	signal cpu_3_data_master_writedata                                       : std_logic_vector(31 downto 0); -- cpu_3:d_writedata -> mm_interconnect_0:cpu_3_data_master_writedata
	signal cpu_4_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_4_data_master_readdata -> cpu_4:d_readdata
	signal cpu_4_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_4_data_master_waitrequest -> cpu_4:d_waitrequest
	signal cpu_4_data_master_debugaccess                                     : std_logic;                     -- cpu_4:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_4_data_master_debugaccess
	signal cpu_4_data_master_address                                         : std_logic_vector(26 downto 0); -- cpu_4:d_address -> mm_interconnect_0:cpu_4_data_master_address
	signal cpu_4_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- cpu_4:d_byteenable -> mm_interconnect_0:cpu_4_data_master_byteenable
	signal cpu_4_data_master_read                                            : std_logic;                     -- cpu_4:d_read -> mm_interconnect_0:cpu_4_data_master_read
	signal cpu_4_data_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:cpu_4_data_master_readdatavalid -> cpu_4:d_readdatavalid
	signal cpu_4_data_master_write                                           : std_logic;                     -- cpu_4:d_write -> mm_interconnect_0:cpu_4_data_master_write
	signal cpu_4_data_master_writedata                                       : std_logic_vector(31 downto 0); -- cpu_4:d_writedata -> mm_interconnect_0:cpu_4_data_master_writedata
	signal cpu_3_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_3_instruction_master_readdata -> cpu_3:i_readdata
	signal cpu_3_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:cpu_3_instruction_master_waitrequest -> cpu_3:i_waitrequest
	signal cpu_3_instruction_master_address                                  : std_logic_vector(26 downto 0); -- cpu_3:i_address -> mm_interconnect_0:cpu_3_instruction_master_address
	signal cpu_3_instruction_master_read                                     : std_logic;                     -- cpu_3:i_read -> mm_interconnect_0:cpu_3_instruction_master_read
	signal cpu_3_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:cpu_3_instruction_master_readdatavalid -> cpu_3:i_readdatavalid
	signal cpu_2_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_2_instruction_master_readdata -> cpu_2:i_readdata
	signal cpu_2_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:cpu_2_instruction_master_waitrequest -> cpu_2:i_waitrequest
	signal cpu_2_instruction_master_address                                  : std_logic_vector(26 downto 0); -- cpu_2:i_address -> mm_interconnect_0:cpu_2_instruction_master_address
	signal cpu_2_instruction_master_read                                     : std_logic;                     -- cpu_2:i_read -> mm_interconnect_0:cpu_2_instruction_master_read
	signal cpu_2_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:cpu_2_instruction_master_readdatavalid -> cpu_2:i_readdatavalid
	signal cpu_1_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_instruction_master_readdata -> cpu_1:i_readdata
	signal cpu_1_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:cpu_1_instruction_master_waitrequest -> cpu_1:i_waitrequest
	signal cpu_1_instruction_master_address                                  : std_logic_vector(26 downto 0); -- cpu_1:i_address -> mm_interconnect_0:cpu_1_instruction_master_address
	signal cpu_1_instruction_master_read                                     : std_logic;                     -- cpu_1:i_read -> mm_interconnect_0:cpu_1_instruction_master_read
	signal cpu_1_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:cpu_1_instruction_master_readdatavalid -> cpu_1:i_readdatavalid
	signal cpu_4_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_4_instruction_master_readdata -> cpu_4:i_readdata
	signal cpu_4_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:cpu_4_instruction_master_waitrequest -> cpu_4:i_waitrequest
	signal cpu_4_instruction_master_address                                  : std_logic_vector(26 downto 0); -- cpu_4:i_address -> mm_interconnect_0:cpu_4_instruction_master_address
	signal cpu_4_instruction_master_read                                     : std_logic;                     -- cpu_4:i_read -> mm_interconnect_0:cpu_4_instruction_master_read
	signal cpu_4_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:cpu_4_instruction_master_readdatavalid -> cpu_4:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect          : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata            : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest         : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write               : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_performance_counter_control_slave_readdata      : std_logic_vector(31 downto 0); -- performance_counter:readdata -> mm_interconnect_0:performance_counter_control_slave_readdata
	signal mm_interconnect_0_performance_counter_control_slave_address       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:performance_counter_control_slave_address -> performance_counter:address
	signal mm_interconnect_0_performance_counter_control_slave_begintransfer : std_logic;                     -- mm_interconnect_0:performance_counter_control_slave_begintransfer -> performance_counter:begintransfer
	signal mm_interconnect_0_performance_counter_control_slave_write         : std_logic;                     -- mm_interconnect_0:performance_counter_control_slave_write -> performance_counter:write
	signal mm_interconnect_0_performance_counter_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:performance_counter_control_slave_writedata -> performance_counter:writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                    : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_1_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- cpu_1:debug_mem_slave_readdata -> mm_interconnect_0:cpu_1_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest               : std_logic;                     -- cpu_1:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_1_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_debugaccess -> cpu_1:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_1_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_address -> cpu_1:debug_mem_slave_address
	signal mm_interconnect_0_cpu_1_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_read -> cpu_1:debug_mem_slave_read
	signal mm_interconnect_0_cpu_1_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_1_debug_mem_slave_byteenable -> cpu_1:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_1_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:cpu_1_debug_mem_slave_write -> cpu_1:debug_mem_slave_write
	signal mm_interconnect_0_cpu_1_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_1_debug_mem_slave_writedata -> cpu_1:debug_mem_slave_writedata
	signal mm_interconnect_0_sdram_controller_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                    : std_logic_vector(15 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest                 : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                     : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                        : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid               : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                       : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                    : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                     : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_mutex_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:mutex_s1_chipselect -> mutex:chipselect
	signal mm_interconnect_0_mutex_s1_readdata                               : std_logic_vector(31 downto 0); -- mutex:data_to_cpu -> mm_interconnect_0:mutex_s1_readdata
	signal mm_interconnect_0_mutex_s1_address                                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:mutex_s1_address -> mutex:address
	signal mm_interconnect_0_mutex_s1_read                                   : std_logic;                     -- mm_interconnect_0:mutex_s1_read -> mutex:read
	signal mm_interconnect_0_mutex_s1_write                                  : std_logic;                     -- mm_interconnect_0:mutex_s1_write -> mutex:write
	signal mm_interconnect_0_mutex_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:mutex_s1_writedata -> mutex:data_from_cpu
	signal mm_interconnect_0_timer1_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:timer1_s1_chipselect -> timer1:chipselect
	signal mm_interconnect_0_timer1_s1_readdata                              : std_logic_vector(15 downto 0); -- timer1:readdata -> mm_interconnect_0:timer1_s1_readdata
	signal mm_interconnect_0_timer1_s1_address                               : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer1_s1_address -> timer1:address
	signal mm_interconnect_0_timer1_s1_write                                 : std_logic;                     -- mm_interconnect_0:timer1_s1_write -> mm_interconnect_0_timer1_s1_write:in
	signal mm_interconnect_0_timer1_s1_writedata                             : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer1_s1_writedata -> timer1:writedata
	signal mm_interconnect_0_cpu_4_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- cpu_4:debug_mem_slave_readdata -> mm_interconnect_0:cpu_4_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_4_debug_mem_slave_waitrequest               : std_logic;                     -- cpu_4:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_4_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_4_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:cpu_4_debug_mem_slave_debugaccess -> cpu_4:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_4_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_4_debug_mem_slave_address -> cpu_4:debug_mem_slave_address
	signal mm_interconnect_0_cpu_4_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:cpu_4_debug_mem_slave_read -> cpu_4:debug_mem_slave_read
	signal mm_interconnect_0_cpu_4_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_4_debug_mem_slave_byteenable -> cpu_4:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_4_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:cpu_4_debug_mem_slave_write -> cpu_4:debug_mem_slave_write
	signal mm_interconnect_0_cpu_4_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_4_debug_mem_slave_writedata -> cpu_4:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_4_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:timer_4_s1_chipselect -> timer_4:chipselect
	signal mm_interconnect_0_timer_4_s1_readdata                             : std_logic_vector(15 downto 0); -- timer_4:readdata -> mm_interconnect_0:timer_4_s1_readdata
	signal mm_interconnect_0_timer_4_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_4_s1_address -> timer_4:address
	signal mm_interconnect_0_timer_4_s1_write                                : std_logic;                     -- mm_interconnect_0:timer_4_s1_write -> mm_interconnect_0_timer_4_s1_write:in
	signal mm_interconnect_0_timer_4_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_4_s1_writedata -> timer_4:writedata
	signal mm_interconnect_0_onchip_memory2_0_s2_chipselect                  : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_chipselect -> onchip_memory2_0:chipselect2
	signal mm_interconnect_0_onchip_memory2_0_s2_readdata                    : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata2 -> mm_interconnect_0:onchip_memory2_0_s2_readdata
	signal mm_interconnect_0_onchip_memory2_0_s2_address                     : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_address -> onchip_memory2_0:address2
	signal mm_interconnect_0_onchip_memory2_0_s2_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s2_byteenable -> onchip_memory2_0:byteenable2
	signal mm_interconnect_0_onchip_memory2_0_s2_write                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_write -> onchip_memory2_0:write2
	signal mm_interconnect_0_onchip_memory2_0_s2_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s2_writedata -> onchip_memory2_0:writedata2
	signal mm_interconnect_0_onchip_memory2_0_s2_clken                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s2_clken -> onchip_memory2_0:clken2
	signal mm_interconnect_0_cpu_3_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- cpu_3:debug_mem_slave_readdata -> mm_interconnect_0:cpu_3_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest               : std_logic;                     -- cpu_3:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_3_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:cpu_3_debug_mem_slave_debugaccess -> cpu_3:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_3_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_3_debug_mem_slave_address -> cpu_3:debug_mem_slave_address
	signal mm_interconnect_0_cpu_3_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:cpu_3_debug_mem_slave_read -> cpu_3:debug_mem_slave_read
	signal mm_interconnect_0_cpu_3_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_3_debug_mem_slave_byteenable -> cpu_3:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_3_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:cpu_3_debug_mem_slave_write -> cpu_3:debug_mem_slave_write
	signal mm_interconnect_0_cpu_3_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_3_debug_mem_slave_writedata -> cpu_3:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_3_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:timer_3_s1_chipselect -> timer_3:chipselect
	signal mm_interconnect_0_timer_3_s1_readdata                             : std_logic_vector(15 downto 0); -- timer_3:readdata -> mm_interconnect_0:timer_3_s1_readdata
	signal mm_interconnect_0_timer_3_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_3_s1_address -> timer_3:address
	signal mm_interconnect_0_timer_3_s1_write                                : std_logic;                     -- mm_interconnect_0:timer_3_s1_write -> mm_interconnect_0_timer_3_s1_write:in
	signal mm_interconnect_0_timer_3_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_3_s1_writedata -> timer_3:writedata
	signal mm_interconnect_0_cpu_2_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- cpu_2:debug_mem_slave_readdata -> mm_interconnect_0:cpu_2_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest               : std_logic;                     -- cpu_2:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_2_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:cpu_2_debug_mem_slave_debugaccess -> cpu_2:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_2_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_2_debug_mem_slave_address -> cpu_2:debug_mem_slave_address
	signal mm_interconnect_0_cpu_2_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:cpu_2_debug_mem_slave_read -> cpu_2:debug_mem_slave_read
	signal mm_interconnect_0_cpu_2_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_2_debug_mem_slave_byteenable -> cpu_2:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_2_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:cpu_2_debug_mem_slave_write -> cpu_2:debug_mem_slave_write
	signal mm_interconnect_0_cpu_2_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_2_debug_mem_slave_writedata -> cpu_2:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_2_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:timer_2_s1_chipselect -> timer_2:chipselect
	signal mm_interconnect_0_timer_2_s1_readdata                             : std_logic_vector(15 downto 0); -- timer_2:readdata -> mm_interconnect_0:timer_2_s1_readdata
	signal mm_interconnect_0_timer_2_s1_address                              : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_2_s1_address -> timer_2:address
	signal mm_interconnect_0_timer_2_s1_write                                : std_logic;                     -- mm_interconnect_0:timer_2_s1_write -> mm_interconnect_0_timer_2_s1_write:in
	signal mm_interconnect_0_timer_2_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_2_s1_writedata -> timer_2:writedata
	signal irq_mapper_receiver0_irq                                          : std_logic;                     -- timer1:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                          : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal cpu_1_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu_1:irq
	signal irq_mapper_001_receiver0_irq                                      : std_logic;                     -- timer_2:irq -> irq_mapper_001:receiver0_irq
	signal cpu_2_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> cpu_2:irq
	signal irq_mapper_002_receiver0_irq                                      : std_logic;                     -- timer_3:irq -> irq_mapper_002:receiver0_irq
	signal cpu_3_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper_002:sender_irq -> cpu_3:irq
	signal irq_mapper_003_receiver0_irq                                      : std_logic;                     -- timer_4:irq -> irq_mapper_003:receiver0_irq
	signal cpu_4_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper_003:sender_irq -> cpu_4:irq
	signal rst_controller_reset_out_reset                                    : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, irq_mapper_001:reset, irq_mapper_002:reset, irq_mapper_003:reset, mm_interconnect_0:cpu_1_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, onchip_memory2_0:reset2, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                : std_logic;                     -- rst_controller:reset_req -> [cpu_1:reset_req, cpu_2:reset_req, cpu_3:reset_req, cpu_4:reset_req, onchip_memory2_0:reset_req, onchip_memory2_0:reset_req2, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                           : std_logic;                     -- reset_reset_n:inv -> [pll:rst, rst_controller:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv     : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv              : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv        : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal mm_interconnect_0_timer1_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_timer1_s1_write:inv -> timer1:write_n
	signal mm_interconnect_0_timer_4_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_timer_4_s1_write:inv -> timer_4:write_n
	signal mm_interconnect_0_timer_3_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_timer_3_s1_write:inv -> timer_3:write_n
	signal mm_interconnect_0_timer_2_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_timer_2_s1_write:inv -> timer_2:write_n
	signal rst_controller_reset_out_reset_ports_inv                          : std_logic;                     -- rst_controller_reset_out_reset:inv -> [cpu_1:reset_n, cpu_2:reset_n, cpu_3:reset_n, cpu_4:reset_n, jtag_uart:rst_n, mutex:reset_n, performance_counter:reset_n, sdram_controller:reset_n, sysid:reset_n, timer1:reset_n, timer_2:reset_n, timer_3:reset_n, timer_4:reset_n]

begin

	cpu_1 : component multicore_cpu_1
		port map (
			clk                                 => pll_outclk0_clk,                                     --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_1_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_1_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_1_data_master_read,                              --                          .read
			d_readdata                          => cpu_1_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_1_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_1_data_master_write,                             --                          .write
			d_writedata                         => cpu_1_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_1_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_1_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_1_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_1_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_1_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_1_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_1_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_1_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_1_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_1_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_1_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_2 : component multicore_cpu_2
		port map (
			clk                                 => pll_outclk0_clk,                                     --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_2_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_2_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_2_data_master_read,                              --                          .read
			d_readdata                          => cpu_2_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_2_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_2_data_master_write,                             --                          .write
			d_writedata                         => cpu_2_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_2_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_2_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_2_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_2_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_2_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_2_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_2_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_2_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_2_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_2_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_2_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_2_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_2_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_2_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_3 : component multicore_cpu_3
		port map (
			clk                                 => pll_outclk0_clk,                                     --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_3_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_3_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_3_data_master_read,                              --                          .read
			d_readdata                          => cpu_3_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_3_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_3_data_master_write,                             --                          .write
			d_writedata                         => cpu_3_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_3_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_3_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_3_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_3_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_3_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_3_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_3_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_3_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_3_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_3_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_3_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_3_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_3_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_3_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	cpu_4 : component multicore_cpu_4
		port map (
			clk                                 => pll_outclk0_clk,                                     --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_4_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_4_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_4_data_master_read,                              --                          .read
			d_readdata                          => cpu_4_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_4_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_4_data_master_write,                             --                          .write
			d_writedata                         => cpu_4_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_4_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_4_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_4_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_4_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_4_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_4_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_4_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_4_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_4_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_4_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_4_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_4_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_4_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_4_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_4_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_4_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	jtag_uart : component multicore_jtag_uart
		port map (
			clk            => pll_outclk0_clk,                                               --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	mutex : component multicore_mutex
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv, -- reset.reset_n
			clk           => pll_outclk0_clk,                          --   clk.clk
			chipselect    => mm_interconnect_0_mutex_s1_chipselect,    --    s1.chipselect
			data_from_cpu => mm_interconnect_0_mutex_s1_writedata,     --      .writedata
			read          => mm_interconnect_0_mutex_s1_read,          --      .read
			write         => mm_interconnect_0_mutex_s1_write,         --      .write
			data_to_cpu   => mm_interconnect_0_mutex_s1_readdata,      --      .readdata
			address       => mm_interconnect_0_mutex_s1_address(0)     --      .address
		);

	onchip_memory2_0 : component multicore_onchip_memory2_0
		port map (
			clk         => pll_outclk0_clk,                                  --   clk1.clk
			address     => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken       => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata    => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,               --       .reset_req
			address2    => mm_interconnect_0_onchip_memory2_0_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_memory2_0_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_memory2_0_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_memory2_0_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_memory2_0_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_memory2_0_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_memory2_0_s2_byteenable, --       .byteenable
			clk2        => pll_outclk0_clk,                                  --   clk2.clk
			reset2      => rst_controller_reset_out_reset,                   -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req                --       .reset_req
		);

	performance_counter : component multicore_performance_counter
		port map (
			clk           => pll_outclk0_clk,                                                   --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                          --         reset.reset_n
			address       => mm_interconnect_0_performance_counter_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_performance_counter_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_performance_counter_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_performance_counter_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_performance_counter_control_slave_writedata      --              .writedata
		);

	pll : component multicore_pll
		port map (
			refclk   => clk_clk,                 --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_outclk0_clk,         -- outclk0.clk
			outclk_1 => sdram_clk_clk,           -- outclk1.clk
			locked   => open                     -- (terminated)
		);

	sdram_controller : component multicore_sdram_controller
		port map (
			clk            => pll_outclk0_clk,                                            --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_wire_addr,                                 --  wire.export
			zs_ba          => sdram_controller_wire_ba,                                   --      .export
			zs_cas_n       => sdram_controller_wire_cas_n,                                --      .export
			zs_cke         => sdram_controller_wire_cke,                                  --      .export
			zs_cs_n        => sdram_controller_wire_cs_n,                                 --      .export
			zs_dq          => sdram_controller_wire_dq,                                   --      .export
			zs_dqm         => sdram_controller_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_controller_wire_ras_n,                                --      .export
			zs_we_n        => sdram_controller_wire_we_n                                  --      .export
		);

	sysid : component multicore_sysid
		port map (
			clock    => pll_outclk0_clk,                                  --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer1 : component multicore_timer1
		port map (
			clk        => pll_outclk0_clk,                             --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    -- reset.reset_n
			address    => mm_interconnect_0_timer1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                     --   irq.irq
		);

	timer_2 : component multicore_timer1
		port map (
			clk        => pll_outclk0_clk,                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_2_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_2_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_2_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_2_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_2_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_001_receiver0_irq                  --   irq.irq
		);

	timer_3 : component multicore_timer1
		port map (
			clk        => pll_outclk0_clk,                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_3_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_3_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_3_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_3_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_3_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_002_receiver0_irq                  --   irq.irq
		);

	timer_4 : component multicore_timer1
		port map (
			clk        => pll_outclk0_clk,                              --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_4_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_4_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_4_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_4_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_4_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_003_receiver0_irq                  --   irq.irq
		);

	mm_interconnect_0 : component multicore_mm_interconnect_0
		port map (
			pll_outclk0_clk                                 => pll_outclk0_clk,                                                   --                       pll_outclk0.clk
			cpu_1_reset_reset_bridge_in_reset_reset         => rst_controller_reset_out_reset,                                    -- cpu_1_reset_reset_bridge_in_reset.reset
			cpu_1_data_master_address                       => cpu_1_data_master_address,                                         --                 cpu_1_data_master.address
			cpu_1_data_master_waitrequest                   => cpu_1_data_master_waitrequest,                                     --                                  .waitrequest
			cpu_1_data_master_byteenable                    => cpu_1_data_master_byteenable,                                      --                                  .byteenable
			cpu_1_data_master_read                          => cpu_1_data_master_read,                                            --                                  .read
			cpu_1_data_master_readdata                      => cpu_1_data_master_readdata,                                        --                                  .readdata
			cpu_1_data_master_readdatavalid                 => cpu_1_data_master_readdatavalid,                                   --                                  .readdatavalid
			cpu_1_data_master_write                         => cpu_1_data_master_write,                                           --                                  .write
			cpu_1_data_master_writedata                     => cpu_1_data_master_writedata,                                       --                                  .writedata
			cpu_1_data_master_debugaccess                   => cpu_1_data_master_debugaccess,                                     --                                  .debugaccess
			cpu_1_instruction_master_address                => cpu_1_instruction_master_address,                                  --          cpu_1_instruction_master.address
			cpu_1_instruction_master_waitrequest            => cpu_1_instruction_master_waitrequest,                              --                                  .waitrequest
			cpu_1_instruction_master_read                   => cpu_1_instruction_master_read,                                     --                                  .read
			cpu_1_instruction_master_readdata               => cpu_1_instruction_master_readdata,                                 --                                  .readdata
			cpu_1_instruction_master_readdatavalid          => cpu_1_instruction_master_readdatavalid,                            --                                  .readdatavalid
			cpu_2_data_master_address                       => cpu_2_data_master_address,                                         --                 cpu_2_data_master.address
			cpu_2_data_master_waitrequest                   => cpu_2_data_master_waitrequest,                                     --                                  .waitrequest
			cpu_2_data_master_byteenable                    => cpu_2_data_master_byteenable,                                      --                                  .byteenable
			cpu_2_data_master_read                          => cpu_2_data_master_read,                                            --                                  .read
			cpu_2_data_master_readdata                      => cpu_2_data_master_readdata,                                        --                                  .readdata
			cpu_2_data_master_readdatavalid                 => cpu_2_data_master_readdatavalid,                                   --                                  .readdatavalid
			cpu_2_data_master_write                         => cpu_2_data_master_write,                                           --                                  .write
			cpu_2_data_master_writedata                     => cpu_2_data_master_writedata,                                       --                                  .writedata
			cpu_2_data_master_debugaccess                   => cpu_2_data_master_debugaccess,                                     --                                  .debugaccess
			cpu_2_instruction_master_address                => cpu_2_instruction_master_address,                                  --          cpu_2_instruction_master.address
			cpu_2_instruction_master_waitrequest            => cpu_2_instruction_master_waitrequest,                              --                                  .waitrequest
			cpu_2_instruction_master_read                   => cpu_2_instruction_master_read,                                     --                                  .read
			cpu_2_instruction_master_readdata               => cpu_2_instruction_master_readdata,                                 --                                  .readdata
			cpu_2_instruction_master_readdatavalid          => cpu_2_instruction_master_readdatavalid,                            --                                  .readdatavalid
			cpu_3_data_master_address                       => cpu_3_data_master_address,                                         --                 cpu_3_data_master.address
			cpu_3_data_master_waitrequest                   => cpu_3_data_master_waitrequest,                                     --                                  .waitrequest
			cpu_3_data_master_byteenable                    => cpu_3_data_master_byteenable,                                      --                                  .byteenable
			cpu_3_data_master_read                          => cpu_3_data_master_read,                                            --                                  .read
			cpu_3_data_master_readdata                      => cpu_3_data_master_readdata,                                        --                                  .readdata
			cpu_3_data_master_readdatavalid                 => cpu_3_data_master_readdatavalid,                                   --                                  .readdatavalid
			cpu_3_data_master_write                         => cpu_3_data_master_write,                                           --                                  .write
			cpu_3_data_master_writedata                     => cpu_3_data_master_writedata,                                       --                                  .writedata
			cpu_3_data_master_debugaccess                   => cpu_3_data_master_debugaccess,                                     --                                  .debugaccess
			cpu_3_instruction_master_address                => cpu_3_instruction_master_address,                                  --          cpu_3_instruction_master.address
			cpu_3_instruction_master_waitrequest            => cpu_3_instruction_master_waitrequest,                              --                                  .waitrequest
			cpu_3_instruction_master_read                   => cpu_3_instruction_master_read,                                     --                                  .read
			cpu_3_instruction_master_readdata               => cpu_3_instruction_master_readdata,                                 --                                  .readdata
			cpu_3_instruction_master_readdatavalid          => cpu_3_instruction_master_readdatavalid,                            --                                  .readdatavalid
			cpu_4_data_master_address                       => cpu_4_data_master_address,                                         --                 cpu_4_data_master.address
			cpu_4_data_master_waitrequest                   => cpu_4_data_master_waitrequest,                                     --                                  .waitrequest
			cpu_4_data_master_byteenable                    => cpu_4_data_master_byteenable,                                      --                                  .byteenable
			cpu_4_data_master_read                          => cpu_4_data_master_read,                                            --                                  .read
			cpu_4_data_master_readdata                      => cpu_4_data_master_readdata,                                        --                                  .readdata
			cpu_4_data_master_readdatavalid                 => cpu_4_data_master_readdatavalid,                                   --                                  .readdatavalid
			cpu_4_data_master_write                         => cpu_4_data_master_write,                                           --                                  .write
			cpu_4_data_master_writedata                     => cpu_4_data_master_writedata,                                       --                                  .writedata
			cpu_4_data_master_debugaccess                   => cpu_4_data_master_debugaccess,                                     --                                  .debugaccess
			cpu_4_instruction_master_address                => cpu_4_instruction_master_address,                                  --          cpu_4_instruction_master.address
			cpu_4_instruction_master_waitrequest            => cpu_4_instruction_master_waitrequest,                              --                                  .waitrequest
			cpu_4_instruction_master_read                   => cpu_4_instruction_master_read,                                     --                                  .read
			cpu_4_instruction_master_readdata               => cpu_4_instruction_master_readdata,                                 --                                  .readdata
			cpu_4_instruction_master_readdatavalid          => cpu_4_instruction_master_readdatavalid,                            --                                  .readdatavalid
			cpu_1_debug_mem_slave_address                   => mm_interconnect_0_cpu_1_debug_mem_slave_address,                   --             cpu_1_debug_mem_slave.address
			cpu_1_debug_mem_slave_write                     => mm_interconnect_0_cpu_1_debug_mem_slave_write,                     --                                  .write
			cpu_1_debug_mem_slave_read                      => mm_interconnect_0_cpu_1_debug_mem_slave_read,                      --                                  .read
			cpu_1_debug_mem_slave_readdata                  => mm_interconnect_0_cpu_1_debug_mem_slave_readdata,                  --                                  .readdata
			cpu_1_debug_mem_slave_writedata                 => mm_interconnect_0_cpu_1_debug_mem_slave_writedata,                 --                                  .writedata
			cpu_1_debug_mem_slave_byteenable                => mm_interconnect_0_cpu_1_debug_mem_slave_byteenable,                --                                  .byteenable
			cpu_1_debug_mem_slave_waitrequest               => mm_interconnect_0_cpu_1_debug_mem_slave_waitrequest,               --                                  .waitrequest
			cpu_1_debug_mem_slave_debugaccess               => mm_interconnect_0_cpu_1_debug_mem_slave_debugaccess,               --                                  .debugaccess
			cpu_2_debug_mem_slave_address                   => mm_interconnect_0_cpu_2_debug_mem_slave_address,                   --             cpu_2_debug_mem_slave.address
			cpu_2_debug_mem_slave_write                     => mm_interconnect_0_cpu_2_debug_mem_slave_write,                     --                                  .write
			cpu_2_debug_mem_slave_read                      => mm_interconnect_0_cpu_2_debug_mem_slave_read,                      --                                  .read
			cpu_2_debug_mem_slave_readdata                  => mm_interconnect_0_cpu_2_debug_mem_slave_readdata,                  --                                  .readdata
			cpu_2_debug_mem_slave_writedata                 => mm_interconnect_0_cpu_2_debug_mem_slave_writedata,                 --                                  .writedata
			cpu_2_debug_mem_slave_byteenable                => mm_interconnect_0_cpu_2_debug_mem_slave_byteenable,                --                                  .byteenable
			cpu_2_debug_mem_slave_waitrequest               => mm_interconnect_0_cpu_2_debug_mem_slave_waitrequest,               --                                  .waitrequest
			cpu_2_debug_mem_slave_debugaccess               => mm_interconnect_0_cpu_2_debug_mem_slave_debugaccess,               --                                  .debugaccess
			cpu_3_debug_mem_slave_address                   => mm_interconnect_0_cpu_3_debug_mem_slave_address,                   --             cpu_3_debug_mem_slave.address
			cpu_3_debug_mem_slave_write                     => mm_interconnect_0_cpu_3_debug_mem_slave_write,                     --                                  .write
			cpu_3_debug_mem_slave_read                      => mm_interconnect_0_cpu_3_debug_mem_slave_read,                      --                                  .read
			cpu_3_debug_mem_slave_readdata                  => mm_interconnect_0_cpu_3_debug_mem_slave_readdata,                  --                                  .readdata
			cpu_3_debug_mem_slave_writedata                 => mm_interconnect_0_cpu_3_debug_mem_slave_writedata,                 --                                  .writedata
			cpu_3_debug_mem_slave_byteenable                => mm_interconnect_0_cpu_3_debug_mem_slave_byteenable,                --                                  .byteenable
			cpu_3_debug_mem_slave_waitrequest               => mm_interconnect_0_cpu_3_debug_mem_slave_waitrequest,               --                                  .waitrequest
			cpu_3_debug_mem_slave_debugaccess               => mm_interconnect_0_cpu_3_debug_mem_slave_debugaccess,               --                                  .debugaccess
			cpu_4_debug_mem_slave_address                   => mm_interconnect_0_cpu_4_debug_mem_slave_address,                   --             cpu_4_debug_mem_slave.address
			cpu_4_debug_mem_slave_write                     => mm_interconnect_0_cpu_4_debug_mem_slave_write,                     --                                  .write
			cpu_4_debug_mem_slave_read                      => mm_interconnect_0_cpu_4_debug_mem_slave_read,                      --                                  .read
			cpu_4_debug_mem_slave_readdata                  => mm_interconnect_0_cpu_4_debug_mem_slave_readdata,                  --                                  .readdata
			cpu_4_debug_mem_slave_writedata                 => mm_interconnect_0_cpu_4_debug_mem_slave_writedata,                 --                                  .writedata
			cpu_4_debug_mem_slave_byteenable                => mm_interconnect_0_cpu_4_debug_mem_slave_byteenable,                --                                  .byteenable
			cpu_4_debug_mem_slave_waitrequest               => mm_interconnect_0_cpu_4_debug_mem_slave_waitrequest,               --                                  .waitrequest
			cpu_4_debug_mem_slave_debugaccess               => mm_interconnect_0_cpu_4_debug_mem_slave_debugaccess,               --                                  .debugaccess
			jtag_uart_avalon_jtag_slave_address             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,             --       jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,               --                                  .write
			jtag_uart_avalon_jtag_slave_read                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                --                                  .read
			jtag_uart_avalon_jtag_slave_readdata            => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,            --                                  .readdata
			jtag_uart_avalon_jtag_slave_writedata           => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,           --                                  .writedata
			jtag_uart_avalon_jtag_slave_waitrequest         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,         --                                  .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect          => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,          --                                  .chipselect
			mutex_s1_address                                => mm_interconnect_0_mutex_s1_address,                                --                          mutex_s1.address
			mutex_s1_write                                  => mm_interconnect_0_mutex_s1_write,                                  --                                  .write
			mutex_s1_read                                   => mm_interconnect_0_mutex_s1_read,                                   --                                  .read
			mutex_s1_readdata                               => mm_interconnect_0_mutex_s1_readdata,                               --                                  .readdata
			mutex_s1_writedata                              => mm_interconnect_0_mutex_s1_writedata,                              --                                  .writedata
			mutex_s1_chipselect                             => mm_interconnect_0_mutex_s1_chipselect,                             --                                  .chipselect
			onchip_memory2_0_s1_address                     => mm_interconnect_0_onchip_memory2_0_s1_address,                     --               onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                       => mm_interconnect_0_onchip_memory2_0_s1_write,                       --                                  .write
			onchip_memory2_0_s1_readdata                    => mm_interconnect_0_onchip_memory2_0_s1_readdata,                    --                                  .readdata
			onchip_memory2_0_s1_writedata                   => mm_interconnect_0_onchip_memory2_0_s1_writedata,                   --                                  .writedata
			onchip_memory2_0_s1_byteenable                  => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                  --                                  .byteenable
			onchip_memory2_0_s1_chipselect                  => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                  --                                  .chipselect
			onchip_memory2_0_s1_clken                       => mm_interconnect_0_onchip_memory2_0_s1_clken,                       --                                  .clken
			onchip_memory2_0_s2_address                     => mm_interconnect_0_onchip_memory2_0_s2_address,                     --               onchip_memory2_0_s2.address
			onchip_memory2_0_s2_write                       => mm_interconnect_0_onchip_memory2_0_s2_write,                       --                                  .write
			onchip_memory2_0_s2_readdata                    => mm_interconnect_0_onchip_memory2_0_s2_readdata,                    --                                  .readdata
			onchip_memory2_0_s2_writedata                   => mm_interconnect_0_onchip_memory2_0_s2_writedata,                   --                                  .writedata
			onchip_memory2_0_s2_byteenable                  => mm_interconnect_0_onchip_memory2_0_s2_byteenable,                  --                                  .byteenable
			onchip_memory2_0_s2_chipselect                  => mm_interconnect_0_onchip_memory2_0_s2_chipselect,                  --                                  .chipselect
			onchip_memory2_0_s2_clken                       => mm_interconnect_0_onchip_memory2_0_s2_clken,                       --                                  .clken
			performance_counter_control_slave_address       => mm_interconnect_0_performance_counter_control_slave_address,       -- performance_counter_control_slave.address
			performance_counter_control_slave_write         => mm_interconnect_0_performance_counter_control_slave_write,         --                                  .write
			performance_counter_control_slave_readdata      => mm_interconnect_0_performance_counter_control_slave_readdata,      --                                  .readdata
			performance_counter_control_slave_writedata     => mm_interconnect_0_performance_counter_control_slave_writedata,     --                                  .writedata
			performance_counter_control_slave_begintransfer => mm_interconnect_0_performance_counter_control_slave_begintransfer, --                                  .begintransfer
			sdram_controller_s1_address                     => mm_interconnect_0_sdram_controller_s1_address,                     --               sdram_controller_s1.address
			sdram_controller_s1_write                       => mm_interconnect_0_sdram_controller_s1_write,                       --                                  .write
			sdram_controller_s1_read                        => mm_interconnect_0_sdram_controller_s1_read,                        --                                  .read
			sdram_controller_s1_readdata                    => mm_interconnect_0_sdram_controller_s1_readdata,                    --                                  .readdata
			sdram_controller_s1_writedata                   => mm_interconnect_0_sdram_controller_s1_writedata,                   --                                  .writedata
			sdram_controller_s1_byteenable                  => mm_interconnect_0_sdram_controller_s1_byteenable,                  --                                  .byteenable
			sdram_controller_s1_readdatavalid               => mm_interconnect_0_sdram_controller_s1_readdatavalid,               --                                  .readdatavalid
			sdram_controller_s1_waitrequest                 => mm_interconnect_0_sdram_controller_s1_waitrequest,                 --                                  .waitrequest
			sdram_controller_s1_chipselect                  => mm_interconnect_0_sdram_controller_s1_chipselect,                  --                                  .chipselect
			sysid_control_slave_address                     => mm_interconnect_0_sysid_control_slave_address,                     --               sysid_control_slave.address
			sysid_control_slave_readdata                    => mm_interconnect_0_sysid_control_slave_readdata,                    --                                  .readdata
			timer1_s1_address                               => mm_interconnect_0_timer1_s1_address,                               --                         timer1_s1.address
			timer1_s1_write                                 => mm_interconnect_0_timer1_s1_write,                                 --                                  .write
			timer1_s1_readdata                              => mm_interconnect_0_timer1_s1_readdata,                              --                                  .readdata
			timer1_s1_writedata                             => mm_interconnect_0_timer1_s1_writedata,                             --                                  .writedata
			timer1_s1_chipselect                            => mm_interconnect_0_timer1_s1_chipselect,                            --                                  .chipselect
			timer_2_s1_address                              => mm_interconnect_0_timer_2_s1_address,                              --                        timer_2_s1.address
			timer_2_s1_write                                => mm_interconnect_0_timer_2_s1_write,                                --                                  .write
			timer_2_s1_readdata                             => mm_interconnect_0_timer_2_s1_readdata,                             --                                  .readdata
			timer_2_s1_writedata                            => mm_interconnect_0_timer_2_s1_writedata,                            --                                  .writedata
			timer_2_s1_chipselect                           => mm_interconnect_0_timer_2_s1_chipselect,                           --                                  .chipselect
			timer_3_s1_address                              => mm_interconnect_0_timer_3_s1_address,                              --                        timer_3_s1.address
			timer_3_s1_write                                => mm_interconnect_0_timer_3_s1_write,                                --                                  .write
			timer_3_s1_readdata                             => mm_interconnect_0_timer_3_s1_readdata,                             --                                  .readdata
			timer_3_s1_writedata                            => mm_interconnect_0_timer_3_s1_writedata,                            --                                  .writedata
			timer_3_s1_chipselect                           => mm_interconnect_0_timer_3_s1_chipselect,                           --                                  .chipselect
			timer_4_s1_address                              => mm_interconnect_0_timer_4_s1_address,                              --                        timer_4_s1.address
			timer_4_s1_write                                => mm_interconnect_0_timer_4_s1_write,                                --                                  .write
			timer_4_s1_readdata                             => mm_interconnect_0_timer_4_s1_readdata,                             --                                  .readdata
			timer_4_s1_writedata                            => mm_interconnect_0_timer_4_s1_writedata,                            --                                  .writedata
			timer_4_s1_chipselect                           => mm_interconnect_0_timer_4_s1_chipselect                            --                                  .chipselect
		);

	irq_mapper : component multicore_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_1_irq_irq                   --    sender.irq
		);

	irq_mapper_001 : component multicore_irq_mapper_001
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq,   -- receiver0.irq
			sender_irq    => cpu_2_irq_irq                   --    sender.irq
		);

	irq_mapper_002 : component multicore_irq_mapper_001
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_002_receiver0_irq,   -- receiver0.irq
			sender_irq    => cpu_3_irq_irq                   --    sender.irq
		);

	irq_mapper_003 : component multicore_irq_mapper_001
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_003_receiver0_irq,   -- receiver0.irq
			sender_irq    => cpu_4_irq_irq                   --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => pll_outclk0_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	mm_interconnect_0_timer1_s1_write_ports_inv <= not mm_interconnect_0_timer1_s1_write;

	mm_interconnect_0_timer_4_s1_write_ports_inv <= not mm_interconnect_0_timer_4_s1_write;

	mm_interconnect_0_timer_3_s1_write_ports_inv <= not mm_interconnect_0_timer_3_s1_write;

	mm_interconnect_0_timer_2_s1_write_ports_inv <= not mm_interconnect_0_timer_2_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of multicore
